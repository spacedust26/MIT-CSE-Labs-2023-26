`timescale 1ns/1ns
`include "csr.v"
module csr_tb;
reg clk,reset;
wire [2:0]w;
csr uut(clk,reset,w);
initial begin
  $dumpfile("csr_tb.vcd");
  $dumpvars(0,csr_tb);
  clk=0;
  forever #10 clk=~clk;
end
initial begin
  reset=1; #20;
  reset=0; #160;
  $display("Test complete");
  $finish;
end
endmodule
